
module crc8_lookup_table (
	input  wire [7:0] address,
	output reg  [7:0] data
);

	always @(*) begin
		case (address)
			8'd000: begin data <= 8'h00; end
			8'd001: begin data <= 8'h07; end
			8'd002: begin data <= 8'h0E; end
			8'd003: begin data <= 8'h09; end
			8'd004: begin data <= 8'h1C; end
			8'd005: begin data <= 8'h1B; end
			8'd006: begin data <= 8'h12; end
			8'd007: begin data <= 8'h15; end
			8'd008: begin data <= 8'h38; end
			8'd009: begin data <= 8'h3F; end
			8'd010: begin data <= 8'h36; end
			8'd011: begin data <= 8'h31; end
			8'd012: begin data <= 8'h24; end
			8'd013: begin data <= 8'h23; end
			8'd014: begin data <= 8'h2A; end
			8'd015: begin data <= 8'h2D; end
			8'd016: begin data <= 8'h70; end
			8'd017: begin data <= 8'h77; end
			8'd018: begin data <= 8'h7E; end
			8'd019: begin data <= 8'h79; end
			8'd020: begin data <= 8'h6C; end
			8'd021: begin data <= 8'h6B; end
			8'd022: begin data <= 8'h62; end
			8'd023: begin data <= 8'h65; end
			8'd024: begin data <= 8'h48; end
			8'd025: begin data <= 8'h4F; end
			8'd026: begin data <= 8'h46; end
			8'd027: begin data <= 8'h41; end
			8'd028: begin data <= 8'h54; end
			8'd029: begin data <= 8'h53; end
			8'd030: begin data <= 8'h5A; end
			8'd031: begin data <= 8'h5D; end
			8'd032: begin data <= 8'hE0; end
			8'd033: begin data <= 8'hE7; end
			8'd034: begin data <= 8'hEE; end
			8'd035: begin data <= 8'hE9; end
			8'd036: begin data <= 8'hFC; end
			8'd037: begin data <= 8'hFB; end
			8'd038: begin data <= 8'hF2; end
			8'd039: begin data <= 8'hF5; end
			8'd040: begin data <= 8'hD8; end
			8'd041: begin data <= 8'hDF; end
			8'd042: begin data <= 8'hD6; end
			8'd043: begin data <= 8'hD1; end
			8'd044: begin data <= 8'hC4; end
			8'd045: begin data <= 8'hC3; end
			8'd046: begin data <= 8'hCA; end
			8'd047: begin data <= 8'hCD; end
			8'd048: begin data <= 8'h90; end
			8'd049: begin data <= 8'h97; end
			8'd050: begin data <= 8'h9E; end
			8'd051: begin data <= 8'h99; end
			8'd052: begin data <= 8'h8C; end
			8'd053: begin data <= 8'h8B; end
			8'd054: begin data <= 8'h82; end
			8'd055: begin data <= 8'h85; end
			8'd056: begin data <= 8'hA8; end
			8'd057: begin data <= 8'hAF; end
			8'd058: begin data <= 8'hA6; end
			8'd059: begin data <= 8'hA1; end
			8'd060: begin data <= 8'hB4; end
			8'd061: begin data <= 8'hB3; end
			8'd062: begin data <= 8'hBA; end
			8'd063: begin data <= 8'hBD; end
			8'd064: begin data <= 8'hC7; end
			8'd065: begin data <= 8'hC0; end
			8'd066: begin data <= 8'hC9; end
			8'd067: begin data <= 8'hCE; end
			8'd068: begin data <= 8'hDB; end
			8'd069: begin data <= 8'hDC; end
			8'd070: begin data <= 8'hD5; end
			8'd071: begin data <= 8'hD2; end
			8'd072: begin data <= 8'hFF; end
			8'd073: begin data <= 8'hF8; end
			8'd074: begin data <= 8'hF1; end
			8'd075: begin data <= 8'hF6; end
			8'd076: begin data <= 8'hE3; end
			8'd077: begin data <= 8'hE4; end
			8'd078: begin data <= 8'hED; end
			8'd079: begin data <= 8'hEA; end
			8'd080: begin data <= 8'hB7; end
			8'd081: begin data <= 8'hB0; end
			8'd082: begin data <= 8'hB9; end
			8'd083: begin data <= 8'hBE; end
			8'd084: begin data <= 8'hAB; end
			8'd085: begin data <= 8'hAC; end
			8'd086: begin data <= 8'hA5; end
			8'd087: begin data <= 8'hA2; end
			8'd088: begin data <= 8'h8F; end
			8'd089: begin data <= 8'h88; end
			8'd090: begin data <= 8'h81; end
			8'd091: begin data <= 8'h86; end
			8'd092: begin data <= 8'h93; end
			8'd093: begin data <= 8'h94; end
			8'd094: begin data <= 8'h9D; end
			8'd095: begin data <= 8'h9A; end
			8'd096: begin data <= 8'h27; end
			8'd097: begin data <= 8'h20; end
			8'd098: begin data <= 8'h29; end
			8'd099: begin data <= 8'h2E; end
			8'd100: begin data <= 8'h3B; end
			8'd101: begin data <= 8'h3C; end
			8'd102: begin data <= 8'h35; end
			8'd103: begin data <= 8'h32; end
			8'd104: begin data <= 8'h1F; end
			8'd105: begin data <= 8'h18; end
			8'd106: begin data <= 8'h11; end
			8'd107: begin data <= 8'h16; end
			8'd108: begin data <= 8'h03; end
			8'd109: begin data <= 8'h04; end
			8'd110: begin data <= 8'h0D; end
			8'd111: begin data <= 8'h0A; end
			8'd112: begin data <= 8'h57; end
			8'd113: begin data <= 8'h50; end
			8'd114: begin data <= 8'h59; end
			8'd115: begin data <= 8'h5E; end
			8'd116: begin data <= 8'h4B; end
			8'd117: begin data <= 8'h4C; end
			8'd118: begin data <= 8'h45; end
			8'd119: begin data <= 8'h42; end
			8'd120: begin data <= 8'h6F; end
			8'd121: begin data <= 8'h68; end
			8'd122: begin data <= 8'h61; end
			8'd123: begin data <= 8'h66; end
			8'd124: begin data <= 8'h73; end
			8'd125: begin data <= 8'h74; end
			8'd126: begin data <= 8'h7D; end
			8'd127: begin data <= 8'h7A; end
			8'd128: begin data <= 8'h89; end
			8'd129: begin data <= 8'h8E; end
			8'd130: begin data <= 8'h87; end
			8'd131: begin data <= 8'h80; end
			8'd132: begin data <= 8'h95; end
			8'd133: begin data <= 8'h92; end
			8'd134: begin data <= 8'h9B; end
			8'd135: begin data <= 8'h9C; end
			8'd136: begin data <= 8'hB1; end
			8'd137: begin data <= 8'hB6; end
			8'd138: begin data <= 8'hBF; end
			8'd139: begin data <= 8'hB8; end
			8'd140: begin data <= 8'hAD; end
			8'd141: begin data <= 8'hAA; end
			8'd142: begin data <= 8'hA3; end
			8'd143: begin data <= 8'hA4; end
			8'd144: begin data <= 8'hF9; end
			8'd145: begin data <= 8'hFE; end
			8'd146: begin data <= 8'hF7; end
			8'd147: begin data <= 8'hF0; end
			8'd148: begin data <= 8'hE5; end
			8'd149: begin data <= 8'hE2; end
			8'd150: begin data <= 8'hEB; end
			8'd151: begin data <= 8'hEC; end
			8'd152: begin data <= 8'hC1; end
			8'd153: begin data <= 8'hC6; end
			8'd154: begin data <= 8'hCF; end
			8'd155: begin data <= 8'hC8; end
			8'd156: begin data <= 8'hDD; end
			8'd157: begin data <= 8'hDA; end
			8'd158: begin data <= 8'hD3; end
			8'd159: begin data <= 8'hD4; end
			8'd160: begin data <= 8'h69; end
			8'd161: begin data <= 8'h6E; end
			8'd162: begin data <= 8'h67; end
			8'd163: begin data <= 8'h60; end
			8'd164: begin data <= 8'h75; end
			8'd165: begin data <= 8'h72; end
			8'd166: begin data <= 8'h7B; end
			8'd167: begin data <= 8'h7C; end
			8'd168: begin data <= 8'h51; end
			8'd169: begin data <= 8'h56; end
			8'd170: begin data <= 8'h5F; end
			8'd171: begin data <= 8'h58; end
			8'd172: begin data <= 8'h4D; end
			8'd173: begin data <= 8'h4A; end
			8'd174: begin data <= 8'h43; end
			8'd175: begin data <= 8'h44; end
			8'd176: begin data <= 8'h19; end
			8'd177: begin data <= 8'h1E; end
			8'd178: begin data <= 8'h17; end
			8'd179: begin data <= 8'h10; end
			8'd180: begin data <= 8'h05; end
			8'd181: begin data <= 8'h02; end
			8'd182: begin data <= 8'h0B; end
			8'd183: begin data <= 8'h0C; end
			8'd184: begin data <= 8'h21; end
			8'd185: begin data <= 8'h26; end
			8'd186: begin data <= 8'h2F; end
			8'd187: begin data <= 8'h28; end
			8'd188: begin data <= 8'h3D; end
			8'd189: begin data <= 8'h3A; end
			8'd190: begin data <= 8'h33; end
			8'd191: begin data <= 8'h34; end
			8'd192: begin data <= 8'h4E; end
			8'd193: begin data <= 8'h49; end
			8'd194: begin data <= 8'h40; end
			8'd195: begin data <= 8'h47; end
			8'd196: begin data <= 8'h52; end
			8'd197: begin data <= 8'h55; end
			8'd198: begin data <= 8'h5C; end
			8'd199: begin data <= 8'h5B; end
			8'd200: begin data <= 8'h76; end
			8'd201: begin data <= 8'h71; end
			8'd202: begin data <= 8'h78; end
			8'd203: begin data <= 8'h7F; end
			8'd204: begin data <= 8'h6A; end
			8'd205: begin data <= 8'h6D; end
			8'd206: begin data <= 8'h64; end
			8'd207: begin data <= 8'h63; end
			8'd208: begin data <= 8'h3E; end
			8'd209: begin data <= 8'h39; end
			8'd210: begin data <= 8'h30; end
			8'd211: begin data <= 8'h37; end
			8'd212: begin data <= 8'h22; end
			8'd213: begin data <= 8'h25; end
			8'd214: begin data <= 8'h2C; end
			8'd215: begin data <= 8'h2B; end
			8'd216: begin data <= 8'h06; end
			8'd217: begin data <= 8'h01; end
			8'd218: begin data <= 8'h08; end
			8'd219: begin data <= 8'h0F; end
			8'd220: begin data <= 8'h1A; end
			8'd221: begin data <= 8'h1D; end
			8'd222: begin data <= 8'h14; end
			8'd223: begin data <= 8'h13; end
			8'd224: begin data <= 8'hAE; end
			8'd225: begin data <= 8'hA9; end
			8'd226: begin data <= 8'hA0; end
			8'd227: begin data <= 8'hA7; end
			8'd228: begin data <= 8'hB2; end
			8'd229: begin data <= 8'hB5; end
			8'd230: begin data <= 8'hBC; end
			8'd231: begin data <= 8'hBB; end
			8'd232: begin data <= 8'h96; end
			8'd233: begin data <= 8'h91; end
			8'd234: begin data <= 8'h98; end
			8'd235: begin data <= 8'h9F; end
			8'd236: begin data <= 8'h8A; end
			8'd237: begin data <= 8'h8D; end
			8'd238: begin data <= 8'h84; end
			8'd239: begin data <= 8'h83; end
			8'd240: begin data <= 8'hDE; end
			8'd241: begin data <= 8'hD9; end
			8'd242: begin data <= 8'hD0; end
			8'd243: begin data <= 8'hD7; end
			8'd244: begin data <= 8'hC2; end
			8'd245: begin data <= 8'hC5; end
			8'd246: begin data <= 8'hCC; end
			8'd247: begin data <= 8'hCB; end
			8'd248: begin data <= 8'hE6; end
			8'd249: begin data <= 8'hE1; end
			8'd250: begin data <= 8'hE8; end
			8'd251: begin data <= 8'hEF; end
			8'd252: begin data <= 8'hFA; end
			8'd253: begin data <= 8'hFD; end
			8'd254: begin data <= 8'hF4; end
			8'd255: begin data <= 8'hF3; end
			
			default: data <= 8'bx;

		endcase
	end

endmodule
