
module crc8_lookup_table (
	input  wire       clk,
	input  wire [7:0] address,
	output reg  [7:0] data
);

	always @(posedge clk) begin
		case (address)
			8'b0000_0000: begin data <= 8'h00; end
			8'b0000_0001: begin data <= 8'h07; end
			8'b0000_0010: begin data <= 8'h0E; end
			8'b0000_0011: begin data <= 8'h09; end
			8'b0000_0100: begin data <= 8'h1C; end
			8'b0000_0101: begin data <= 8'h1B; end
			8'b0000_0110: begin data <= 8'h12; end
			8'b0000_0111: begin data <= 8'h15; end
			8'b0000_1000: begin data <= 8'h38; end
			8'b0000_1001: begin data <= 8'h3F; end
			8'b0000_1010: begin data <= 8'h36; end
			8'b0000_1011: begin data <= 8'h31; end
			8'b0000_1100: begin data <= 8'h24; end
			8'b0000_1101: begin data <= 8'h23; end
			8'b0000_1110: begin data <= 8'h2A; end
			8'b0000_1111: begin data <= 8'h2D; end
			8'b0001_0000: begin data <= 8'h70; end
			8'b0001_0001: begin data <= 8'h77; end
			8'b0001_0010: begin data <= 8'h7E; end
			8'b0001_0011: begin data <= 8'h79; end
			8'b0001_0100: begin data <= 8'h6C; end
			8'b0001_0101: begin data <= 8'h6B; end
			8'b0001_0110: begin data <= 8'h62; end
			8'b0001_0111: begin data <= 8'h65; end
			8'b0001_1000: begin data <= 8'h48; end
			8'b0001_1001: begin data <= 8'h4F; end
			8'b0001_1010: begin data <= 8'h46; end
			8'b0001_1011: begin data <= 8'h41; end
			8'b0001_1100: begin data <= 8'h54; end
			8'b0001_1101: begin data <= 8'h53; end
			8'b0001_1110: begin data <= 8'h5A; end
			8'b0001_1111: begin data <= 8'h5D; end
			8'b0010_0000: begin data <= 8'hE0; end
			8'b0010_0001: begin data <= 8'hE7; end
			8'b0010_0010: begin data <= 8'hEE; end
			8'b0010_0011: begin data <= 8'hE9; end
			8'b0010_0100: begin data <= 8'hFC; end
			8'b0010_0101: begin data <= 8'hFB; end
			8'b0010_0110: begin data <= 8'hF2; end
			8'b0010_0111: begin data <= 8'hF5; end
			8'b0010_1000: begin data <= 8'hD8; end
			8'b0010_1001: begin data <= 8'hDF; end
			8'b0010_1010: begin data <= 8'hD6; end
			8'b0010_1011: begin data <= 8'hD1; end
			8'b0010_1100: begin data <= 8'hC4; end
			8'b0010_1101: begin data <= 8'hC3; end
			8'b0010_1110: begin data <= 8'hCA; end
			8'b0010_1111: begin data <= 8'hCD; end
			8'b0011_0000: begin data <= 8'h90; end
			8'b0011_0001: begin data <= 8'h97; end
			8'b0011_0010: begin data <= 8'h9E; end
			8'b0011_0011: begin data <= 8'h99; end
			8'b0011_0100: begin data <= 8'h8C; end
			8'b0011_0101: begin data <= 8'h8B; end
			8'b0011_0110: begin data <= 8'h82; end
			8'b0011_0111: begin data <= 8'h85; end
			8'b0011_1000: begin data <= 8'hA8; end
			8'b0011_1001: begin data <= 8'hAF; end
			8'b0011_1010: begin data <= 8'hA6; end
			8'b0011_1011: begin data <= 8'hA1; end
			8'b0011_1100: begin data <= 8'hB4; end
			8'b0011_1101: begin data <= 8'hB3; end
			8'b0011_1110: begin data <= 8'hBA; end
			8'b0011_1111: begin data <= 8'hBD; end
			8'b0100_0000: begin data <= 8'hC7; end
			8'b0100_0001: begin data <= 8'hC0; end
			8'b0100_0010: begin data <= 8'hC9; end
			8'b0100_0011: begin data <= 8'hCE; end
			8'b0100_0100: begin data <= 8'hDB; end
			8'b0100_0101: begin data <= 8'hDC; end
			8'b0100_0110: begin data <= 8'hD5; end
			8'b0100_0111: begin data <= 8'hD2; end
			8'b0100_1000: begin data <= 8'hFF; end
			8'b0100_1001: begin data <= 8'hF8; end
			8'b0100_1010: begin data <= 8'hF1; end
			8'b0100_1011: begin data <= 8'hF6; end
			8'b0100_1100: begin data <= 8'hE3; end
			8'b0100_1101: begin data <= 8'hE4; end
			8'b0100_1110: begin data <= 8'hED; end
			8'b0100_1111: begin data <= 8'hEA; end
			8'b0101_0000: begin data <= 8'hB7; end
			8'b0101_0001: begin data <= 8'hB0; end
			8'b0101_0010: begin data <= 8'hB9; end
			8'b0101_0011: begin data <= 8'hBE; end
			8'b0101_0100: begin data <= 8'hAB; end
			8'b0101_0101: begin data <= 8'hAC; end
			8'b0101_0110: begin data <= 8'hA5; end
			8'b0101_0111: begin data <= 8'hA2; end
			8'b0101_1000: begin data <= 8'h8F; end
			8'b0101_1001: begin data <= 8'h88; end
			8'b0101_1010: begin data <= 8'h81; end
			8'b0101_1011: begin data <= 8'h86; end
			8'b0101_1100: begin data <= 8'h93; end
			8'b0101_1101: begin data <= 8'h94; end
			8'b0101_1110: begin data <= 8'h9D; end
			8'b0101_1111: begin data <= 8'h9A; end
			8'b0110_0000: begin data <= 8'h27; end
			8'b0110_0001: begin data <= 8'h20; end
			8'b0110_0010: begin data <= 8'h29; end
			8'b0110_0011: begin data <= 8'h2E; end
			8'b0110_0100: begin data <= 8'h3B; end
			8'b0110_0101: begin data <= 8'h3C; end
			8'b0110_0110: begin data <= 8'h35; end
			8'b0110_0111: begin data <= 8'h32; end
			8'b0110_1000: begin data <= 8'h1F; end
			8'b0110_1001: begin data <= 8'h18; end
			8'b0110_1010: begin data <= 8'h11; end
			8'b0110_1011: begin data <= 8'h16; end
			8'b0110_1100: begin data <= 8'h03; end
			8'b0110_1101: begin data <= 8'h04; end
			8'b0110_1110: begin data <= 8'h0D; end
			8'b0110_1111: begin data <= 8'h0A; end
			8'b0111_0000: begin data <= 8'h57; end
			8'b0111_0001: begin data <= 8'h50; end
			8'b0111_0010: begin data <= 8'h59; end
			8'b0111_0011: begin data <= 8'h5E; end
			8'b0111_0100: begin data <= 8'h4B; end
			8'b0111_0101: begin data <= 8'h4C; end
			8'b0111_0110: begin data <= 8'h45; end
			8'b0111_0111: begin data <= 8'h42; end
			8'b0111_1000: begin data <= 8'h6F; end
			8'b0111_1001: begin data <= 8'h68; end
			8'b0111_1010: begin data <= 8'h61; end
			8'b0111_1011: begin data <= 8'h66; end
			8'b0111_1100: begin data <= 8'h73; end
			8'b0111_1101: begin data <= 8'h74; end
			8'b0111_1110: begin data <= 8'h7D; end
			8'b0111_1111: begin data <= 8'h7A; end
			8'b1000_0000: begin data <= 8'h89; end
			8'b1000_0001: begin data <= 8'h8E; end
			8'b1000_0010: begin data <= 8'h87; end
			8'b1000_0011: begin data <= 8'h80; end
			8'b1000_0100: begin data <= 8'h95; end
			8'b1000_0101: begin data <= 8'h92; end
			8'b1000_0110: begin data <= 8'h9B; end
			8'b1000_0111: begin data <= 8'h9C; end
			8'b1000_1000: begin data <= 8'hB1; end
			8'b1000_1001: begin data <= 8'hB6; end
			8'b1000_1010: begin data <= 8'hBF; end
			8'b1000_1011: begin data <= 8'hB8; end
			8'b1000_1100: begin data <= 8'hAD; end
			8'b1000_1101: begin data <= 8'hAA; end
			8'b1000_1110: begin data <= 8'hA3; end
			8'b1000_1111: begin data <= 8'hA4; end
			8'b1001_0000: begin data <= 8'hF9; end
			8'b1001_0001: begin data <= 8'hFE; end
			8'b1001_0010: begin data <= 8'hF7; end
			8'b1001_0011: begin data <= 8'hF0; end
			8'b1001_0100: begin data <= 8'hE5; end
			8'b1001_0101: begin data <= 8'hE2; end
			8'b1001_0110: begin data <= 8'hEB; end
			8'b1001_0111: begin data <= 8'hEC; end
			8'b1001_1000: begin data <= 8'hC1; end
			8'b1001_1001: begin data <= 8'hC6; end
			8'b1001_1010: begin data <= 8'hCF; end
			8'b1001_1011: begin data <= 8'hC8; end
			8'b1001_1100: begin data <= 8'hDD; end
			8'b1001_1101: begin data <= 8'hDA; end
			8'b1001_1110: begin data <= 8'hD3; end
			8'b1001_1111: begin data <= 8'hD4; end
			8'b1010_0000: begin data <= 8'h69; end
			8'b1010_0001: begin data <= 8'h6E; end
			8'b1010_0010: begin data <= 8'h67; end
			8'b1010_0011: begin data <= 8'h60; end
			8'b1010_0100: begin data <= 8'h75; end
			8'b1010_0101: begin data <= 8'h72; end
			8'b1010_0110: begin data <= 8'h7B; end
			8'b1010_0111: begin data <= 8'h7C; end
			8'b1010_1000: begin data <= 8'h51; end
			8'b1010_1001: begin data <= 8'h56; end
			8'b1010_1010: begin data <= 8'h5F; end
			8'b1010_1011: begin data <= 8'h58; end
			8'b1010_1100: begin data <= 8'h4D; end
			8'b1010_1101: begin data <= 8'h4A; end
			8'b1010_1110: begin data <= 8'h43; end
			8'b1010_1111: begin data <= 8'h44; end
			8'b1011_0000: begin data <= 8'h19; end
			8'b1011_0001: begin data <= 8'h1E; end
			8'b1011_0010: begin data <= 8'h17; end
			8'b1011_0011: begin data <= 8'h10; end
			8'b1011_0100: begin data <= 8'h05; end
			8'b1011_0101: begin data <= 8'h02; end
			8'b1011_0110: begin data <= 8'h0B; end
			8'b1011_0111: begin data <= 8'h0C; end
			8'b1011_1000: begin data <= 8'h21; end
			8'b1011_1001: begin data <= 8'h26; end
			8'b1011_1010: begin data <= 8'h2F; end
			8'b1011_1011: begin data <= 8'h28; end
			8'b1011_1100: begin data <= 8'h3D; end
			8'b1011_1101: begin data <= 8'h3A; end
			8'b1011_1110: begin data <= 8'h33; end
			8'b1011_1111: begin data <= 8'h34; end
			8'b1100_0000: begin data <= 8'h4E; end
			8'b1100_0001: begin data <= 8'h49; end
			8'b1100_0010: begin data <= 8'h40; end
			8'b1100_0011: begin data <= 8'h47; end
			8'b1100_0100: begin data <= 8'h52; end
			8'b1100_0101: begin data <= 8'h55; end
			8'b1100_0110: begin data <= 8'h5C; end
			8'b1100_0111: begin data <= 8'h5B; end
			8'b1100_1000: begin data <= 8'h76; end
			8'b1100_1001: begin data <= 8'h71; end
			8'b1100_1010: begin data <= 8'h78; end
			8'b1100_1011: begin data <= 8'h7F; end
			8'b1100_1100: begin data <= 8'h6A; end
			8'b1100_1101: begin data <= 8'h6D; end
			8'b1100_1110: begin data <= 8'h64; end
			8'b1100_1111: begin data <= 8'h63; end
			8'b1101_0000: begin data <= 8'h3E; end
			8'b1101_0001: begin data <= 8'h39; end
			8'b1101_0010: begin data <= 8'h30; end
			8'b1101_0011: begin data <= 8'h37; end
			8'b1101_0100: begin data <= 8'h22; end
			8'b1101_0101: begin data <= 8'h25; end
			8'b1101_0110: begin data <= 8'h2C; end
			8'b1101_0111: begin data <= 8'h2B; end
			8'b1101_1000: begin data <= 8'h06; end
			8'b1101_1001: begin data <= 8'h01; end
			8'b1101_1010: begin data <= 8'h08; end
			8'b1101_1011: begin data <= 8'h0F; end
			8'b1101_1100: begin data <= 8'h1A; end
			8'b1101_1101: begin data <= 8'h1D; end
			8'b1101_1110: begin data <= 8'h14; end
			8'b1101_1111: begin data <= 8'h13; end
			8'b1110_0000: begin data <= 8'hAE; end
			8'b1110_0001: begin data <= 8'hA9; end
			8'b1110_0010: begin data <= 8'hA0; end
			8'b1110_0011: begin data <= 8'hA7; end
			8'b1110_0100: begin data <= 8'hB2; end
			8'b1110_0101: begin data <= 8'hB5; end
			8'b1110_0110: begin data <= 8'hBC; end
			8'b1110_0111: begin data <= 8'hBB; end
			8'b1110_1000: begin data <= 8'h96; end
			8'b1110_1001: begin data <= 8'h91; end
			8'b1110_1010: begin data <= 8'h98; end
			8'b1110_1011: begin data <= 8'h9F; end
			8'b1110_1100: begin data <= 8'h8A; end
			8'b1110_1101: begin data <= 8'h8D; end
			8'b1110_1110: begin data <= 8'h84; end
			8'b1110_1111: begin data <= 8'h83; end
			8'b1111_0000: begin data <= 8'hDE; end
			8'b1111_0001: begin data <= 8'hD9; end
			8'b1111_0010: begin data <= 8'hD0; end
			8'b1111_0011: begin data <= 8'hD7; end
			8'b1111_0100: begin data <= 8'hC2; end
			8'b1111_0101: begin data <= 8'hC5; end
			8'b1111_0110: begin data <= 8'hCC; end
			8'b1111_0111: begin data <= 8'hCB; end
			8'b1111_1000: begin data <= 8'hE6; end
			8'b1111_1001: begin data <= 8'hE1; end
			8'b1111_1010: begin data <= 8'hE8; end
			8'b1111_1011: begin data <= 8'hEF; end
			8'b1111_1100: begin data <= 8'hFA; end
			8'b1111_1101: begin data <= 8'hFD; end
			8'b1111_1110: begin data <= 8'hF4; end
			8'b1111_1111: begin data <= 8'hF3; end
			
			default: data <= 8'bx;
		endcase
	end

endmodule
