
module encoder_8b10b_rom (

	input  wire [7:0] data_in,
	input  wire       current_rd,
	input  wire       KI,
	output reg  [9:0] code,
	output reg        next_rd

);

	parameter same = 1'b0;
	parameter flip = 1'b1;

	always @(*) begin
		case ({data_in, current_rd, KI})
			10'b000_00000_0_0: begin code = 10'b100111_0100; next_rd = same; end
			10'b000_00000_1_0: begin code = 10'b011000_1011; next_rd = same; end
			10'b001_00000_0_0: begin code = 10'b100111_1001; next_rd = flip; end
			10'b001_00000_1_0: begin code = 10'b011000_1001; next_rd = flip; end
			10'b010_00000_0_0: begin code = 10'b100111_0101; next_rd = flip; end
			10'b010_00000_1_0: begin code = 10'b011000_0101; next_rd = flip; end
			10'b011_00000_0_0: begin code = 10'b100111_0011; next_rd = flip; end
			10'b011_00000_1_0: begin code = 10'b011000_1100; next_rd = flip; end
			10'b100_00000_0_0: begin code = 10'b100111_0010; next_rd = same; end
			10'b100_00000_1_0: begin code = 10'b011000_1101; next_rd = same; end
			10'b101_00000_0_0: begin code = 10'b100111_1010; next_rd = flip; end
			10'b101_00000_1_0: begin code = 10'b011000_1010; next_rd = flip; end
			10'b110_00000_0_0: begin code = 10'b100111_0110; next_rd = flip; end
			10'b110_00000_1_0: begin code = 10'b011000_0110; next_rd = flip; end
			10'b111_00000_0_0: begin code = 10'b100111_0001; next_rd = same; end
			10'b111_00000_1_0: begin code = 10'b011000_1110; next_rd = same; end
			10'b000_00001_0_0: begin code = 10'b011101_0100; next_rd = same; end
			10'b000_00001_1_0: begin code = 10'b100010_1011; next_rd = same; end
			10'b001_00001_0_0: begin code = 10'b011101_1001; next_rd = flip; end
			10'b001_00001_1_0: begin code = 10'b100010_1001; next_rd = flip; end
			10'b010_00001_0_0: begin code = 10'b011101_0101; next_rd = flip; end
			10'b010_00001_1_0: begin code = 10'b100010_0101; next_rd = flip; end
			10'b011_00001_0_0: begin code = 10'b011101_0011; next_rd = flip; end
			10'b011_00001_1_0: begin code = 10'b100010_1100; next_rd = flip; end
			10'b100_00001_0_0: begin code = 10'b011101_0010; next_rd = same; end
			10'b100_00001_1_0: begin code = 10'b100010_1101; next_rd = same; end
			10'b101_00001_0_0: begin code = 10'b011101_1010; next_rd = flip; end
			10'b101_00001_1_0: begin code = 10'b100010_1010; next_rd = flip; end
			10'b110_00001_0_0: begin code = 10'b011101_0110; next_rd = flip; end
			10'b110_00001_1_0: begin code = 10'b100010_0110; next_rd = flip; end
			10'b111_00001_0_0: begin code = 10'b011101_0001; next_rd = same; end
			10'b111_00001_1_0: begin code = 10'b100010_1110; next_rd = same; end
			10'b000_00010_0_0: begin code = 10'b101101_0100; next_rd = same; end
			10'b000_00010_1_0: begin code = 10'b010010_1011; next_rd = same; end
			10'b001_00010_0_0: begin code = 10'b101101_1001; next_rd = flip; end
			10'b001_00010_1_0: begin code = 10'b010010_1001; next_rd = flip; end
			10'b010_00010_0_0: begin code = 10'b101101_0101; next_rd = flip; end
			10'b010_00010_1_0: begin code = 10'b010010_0101; next_rd = flip; end
			10'b011_00010_0_0: begin code = 10'b101101_0011; next_rd = flip; end
			10'b011_00010_1_0: begin code = 10'b010010_1100; next_rd = flip; end
			10'b100_00010_0_0: begin code = 10'b101101_0010; next_rd = same; end
			10'b100_00010_1_0: begin code = 10'b010010_1101; next_rd = same; end
			10'b101_00010_0_0: begin code = 10'b101101_1010; next_rd = flip; end
			10'b101_00010_1_0: begin code = 10'b010010_1010; next_rd = flip; end
			10'b110_00010_0_0: begin code = 10'b101101_0110; next_rd = flip; end
			10'b110_00010_1_0: begin code = 10'b010010_0110; next_rd = flip; end
			10'b111_00010_0_0: begin code = 10'b101101_0001; next_rd = same; end
			10'b111_00010_1_0: begin code = 10'b010010_1110; next_rd = same; end
			10'b000_00011_0_0: begin code = 10'b110001_1011; next_rd = flip; end
			10'b000_00011_1_0: begin code = 10'b110001_0100; next_rd = flip; end
			10'b001_00011_0_0: begin code = 10'b110001_1001; next_rd = same; end
			10'b001_00011_1_0: begin code = 10'b110001_1001; next_rd = same; end
			10'b010_00011_0_0: begin code = 10'b110001_0101; next_rd = same; end
			10'b010_00011_1_0: begin code = 10'b110001_0101; next_rd = same; end
			10'b011_00011_0_0: begin code = 10'b110001_1100; next_rd = same; end
			10'b011_00011_1_0: begin code = 10'b110001_0011; next_rd = same; end
			10'b100_00011_0_0: begin code = 10'b110001_1101; next_rd = flip; end
			10'b100_00011_1_0: begin code = 10'b110001_0010; next_rd = flip; end
			10'b101_00011_0_0: begin code = 10'b110001_1010; next_rd = same; end
			10'b101_00011_1_0: begin code = 10'b110001_1010; next_rd = same; end
			10'b110_00011_0_0: begin code = 10'b110001_0110; next_rd = same; end
			10'b110_00011_1_0: begin code = 10'b110001_0110; next_rd = same; end
			10'b111_00011_0_0: begin code = 10'b110001_1110; next_rd = flip; end
			10'b111_00011_1_0: begin code = 10'b110001_0001; next_rd = flip; end
			10'b000_00100_0_0: begin code = 10'b110101_0100; next_rd = same; end
			10'b000_00100_1_0: begin code = 10'b001010_1011; next_rd = same; end
			10'b001_00100_0_0: begin code = 10'b110101_1001; next_rd = flip; end
			10'b001_00100_1_0: begin code = 10'b001010_1001; next_rd = flip; end
			10'b010_00100_0_0: begin code = 10'b110101_0101; next_rd = flip; end
			10'b010_00100_1_0: begin code = 10'b001010_0101; next_rd = flip; end
			10'b011_00100_0_0: begin code = 10'b110101_0011; next_rd = flip; end
			10'b011_00100_1_0: begin code = 10'b001010_1100; next_rd = flip; end
			10'b100_00100_0_0: begin code = 10'b110101_0010; next_rd = same; end
			10'b100_00100_1_0: begin code = 10'b001010_1101; next_rd = same; end
			10'b101_00100_0_0: begin code = 10'b110101_1010; next_rd = flip; end
			10'b101_00100_1_0: begin code = 10'b001010_1010; next_rd = flip; end
			10'b110_00100_0_0: begin code = 10'b110101_0110; next_rd = flip; end
			10'b110_00100_1_0: begin code = 10'b001010_0110; next_rd = flip; end
			10'b111_00100_0_0: begin code = 10'b110101_0001; next_rd = same; end
			10'b111_00100_1_0: begin code = 10'b001010_1110; next_rd = same; end
			10'b000_00101_0_0: begin code = 10'b101001_1011; next_rd = flip; end
			10'b000_00101_1_0: begin code = 10'b101001_0100; next_rd = flip; end
			10'b001_00101_0_0: begin code = 10'b101001_1001; next_rd = same; end
			10'b001_00101_1_0: begin code = 10'b101001_1001; next_rd = same; end
			10'b010_00101_0_0: begin code = 10'b101001_0101; next_rd = same; end
			10'b010_00101_1_0: begin code = 10'b101001_0101; next_rd = same; end
			10'b011_00101_0_0: begin code = 10'b101001_1100; next_rd = same; end
			10'b011_00101_1_0: begin code = 10'b101001_0011; next_rd = same; end
			10'b100_00101_0_0: begin code = 10'b101001_1101; next_rd = flip; end
			10'b100_00101_1_0: begin code = 10'b101001_0010; next_rd = flip; end
			10'b101_00101_0_0: begin code = 10'b101001_1010; next_rd = same; end
			10'b101_00101_1_0: begin code = 10'b101001_1010; next_rd = same; end
			10'b110_00101_0_0: begin code = 10'b101001_0110; next_rd = same; end
			10'b110_00101_1_0: begin code = 10'b101001_0110; next_rd = same; end
			10'b111_00101_0_0: begin code = 10'b101001_1110; next_rd = flip; end
			10'b111_00101_1_0: begin code = 10'b101001_0001; next_rd = flip; end
			10'b000_00110_0_0: begin code = 10'b011001_1011; next_rd = flip; end
			10'b000_00110_1_0: begin code = 10'b011001_0100; next_rd = flip; end
			10'b001_00110_0_0: begin code = 10'b011001_1001; next_rd = same; end
			10'b001_00110_1_0: begin code = 10'b011001_1001; next_rd = same; end
			10'b010_00110_0_0: begin code = 10'b011001_0101; next_rd = same; end
			10'b010_00110_1_0: begin code = 10'b011001_0101; next_rd = same; end
			10'b011_00110_0_0: begin code = 10'b011001_1100; next_rd = same; end
			10'b011_00110_1_0: begin code = 10'b011001_0011; next_rd = same; end
			10'b100_00110_0_0: begin code = 10'b011001_1101; next_rd = flip; end
			10'b100_00110_1_0: begin code = 10'b011001_0010; next_rd = flip; end
			10'b101_00110_0_0: begin code = 10'b011001_1010; next_rd = same; end
			10'b101_00110_1_0: begin code = 10'b011001_1010; next_rd = same; end
			10'b110_00110_0_0: begin code = 10'b011001_0110; next_rd = same; end
			10'b110_00110_1_0: begin code = 10'b011001_0110; next_rd = same; end
			10'b111_00110_0_0: begin code = 10'b011001_1110; next_rd = flip; end
			10'b111_00110_1_0: begin code = 10'b011001_0001; next_rd = flip; end
			10'b000_00111_0_0: begin code = 10'b111000_1011; next_rd = flip; end
			10'b000_00111_1_0: begin code = 10'b000111_0100; next_rd = flip; end
			10'b001_00111_0_0: begin code = 10'b111000_1001; next_rd = same; end
			10'b001_00111_1_0: begin code = 10'b000111_1001; next_rd = same; end
			10'b010_00111_0_0: begin code = 10'b111000_0101; next_rd = same; end
			10'b010_00111_1_0: begin code = 10'b000111_0101; next_rd = same; end
			10'b011_00111_0_0: begin code = 10'b111000_1100; next_rd = same; end
			10'b011_00111_1_0: begin code = 10'b000111_0011; next_rd = same; end
			10'b100_00111_0_0: begin code = 10'b111000_1101; next_rd = flip; end
			10'b100_00111_1_0: begin code = 10'b000111_0010; next_rd = flip; end
			10'b101_00111_0_0: begin code = 10'b111000_1010; next_rd = same; end
			10'b101_00111_1_0: begin code = 10'b000111_1010; next_rd = same; end
			10'b110_00111_0_0: begin code = 10'b111000_0110; next_rd = same; end
			10'b110_00111_1_0: begin code = 10'b000111_0110; next_rd = same; end
			10'b111_00111_0_0: begin code = 10'b111000_1110; next_rd = flip; end
			10'b111_00111_1_0: begin code = 10'b000111_0001; next_rd = flip; end
			10'b000_01000_0_0: begin code = 10'b111001_0100; next_rd = same; end
			10'b000_01000_1_0: begin code = 10'b000110_1011; next_rd = same; end
			10'b001_01000_0_0: begin code = 10'b111001_1001; next_rd = flip; end
			10'b001_01000_1_0: begin code = 10'b000110_1001; next_rd = flip; end
			10'b010_01000_0_0: begin code = 10'b111001_0101; next_rd = flip; end
			10'b010_01000_1_0: begin code = 10'b000110_0101; next_rd = flip; end
			10'b011_01000_0_0: begin code = 10'b111001_0011; next_rd = flip; end
			10'b011_01000_1_0: begin code = 10'b000110_1100; next_rd = flip; end
			10'b100_01000_0_0: begin code = 10'b111001_0010; next_rd = same; end
			10'b100_01000_1_0: begin code = 10'b000110_1101; next_rd = same; end
			10'b101_01000_0_0: begin code = 10'b111001_1010; next_rd = flip; end
			10'b101_01000_1_0: begin code = 10'b000110_1010; next_rd = flip; end
			10'b110_01000_0_0: begin code = 10'b111001_0110; next_rd = flip; end
			10'b110_01000_1_0: begin code = 10'b000110_0110; next_rd = flip; end
			10'b111_01000_0_0: begin code = 10'b111001_0001; next_rd = same; end
			10'b111_01000_1_0: begin code = 10'b000110_1110; next_rd = same; end
			10'b000_01001_0_0: begin code = 10'b100101_1011; next_rd = flip; end
			10'b000_01001_1_0: begin code = 10'b100101_0100; next_rd = flip; end
			10'b001_01001_0_0: begin code = 10'b100101_1001; next_rd = same; end
			10'b001_01001_1_0: begin code = 10'b100101_1001; next_rd = same; end
			10'b010_01001_0_0: begin code = 10'b100101_0101; next_rd = same; end
			10'b010_01001_1_0: begin code = 10'b100101_0101; next_rd = same; end
			10'b011_01001_0_0: begin code = 10'b100101_1100; next_rd = same; end
			10'b011_01001_1_0: begin code = 10'b100101_0011; next_rd = same; end
			10'b100_01001_0_0: begin code = 10'b100101_1101; next_rd = flip; end
			10'b100_01001_1_0: begin code = 10'b100101_0010; next_rd = flip; end
			10'b101_01001_0_0: begin code = 10'b100101_1010; next_rd = same; end
			10'b101_01001_1_0: begin code = 10'b100101_1010; next_rd = same; end
			10'b110_01001_0_0: begin code = 10'b100101_0110; next_rd = same; end
			10'b110_01001_1_0: begin code = 10'b100101_0110; next_rd = same; end
			10'b111_01001_0_0: begin code = 10'b100101_1110; next_rd = flip; end
			10'b111_01001_1_0: begin code = 10'b100101_0001; next_rd = flip; end
			10'b000_01010_0_0: begin code = 10'b010101_1011; next_rd = flip; end
			10'b000_01010_1_0: begin code = 10'b010101_0100; next_rd = flip; end
			10'b001_01010_0_0: begin code = 10'b010101_1001; next_rd = same; end
			10'b001_01010_1_0: begin code = 10'b010101_1001; next_rd = same; end
			10'b010_01010_0_0: begin code = 10'b010101_0101; next_rd = same; end
			10'b010_01010_1_0: begin code = 10'b010101_0101; next_rd = same; end
			10'b011_01010_0_0: begin code = 10'b010101_1100; next_rd = same; end
			10'b011_01010_1_0: begin code = 10'b010101_0011; next_rd = same; end
			10'b100_01010_0_0: begin code = 10'b010101_1101; next_rd = flip; end
			10'b100_01010_1_0: begin code = 10'b010101_0010; next_rd = flip; end
			10'b101_01010_0_0: begin code = 10'b010101_1010; next_rd = same; end
			10'b101_01010_1_0: begin code = 10'b010101_1010; next_rd = same; end
			10'b110_01010_0_0: begin code = 10'b010101_0110; next_rd = same; end
			10'b110_01010_1_0: begin code = 10'b010101_0110; next_rd = same; end
			10'b111_01010_0_0: begin code = 10'b010101_1110; next_rd = flip; end
			10'b111_01010_1_0: begin code = 10'b010101_0001; next_rd = flip; end
			10'b000_01011_0_0: begin code = 10'b110100_1011; next_rd = flip; end
			10'b000_01011_1_0: begin code = 10'b110100_0100; next_rd = flip; end
			10'b001_01011_0_0: begin code = 10'b110100_1001; next_rd = same; end
			10'b001_01011_1_0: begin code = 10'b110100_1001; next_rd = same; end
			10'b010_01011_0_0: begin code = 10'b110100_0101; next_rd = same; end
			10'b010_01011_1_0: begin code = 10'b110100_0101; next_rd = same; end
			10'b011_01011_0_0: begin code = 10'b110100_1100; next_rd = same; end
			10'b011_01011_1_0: begin code = 10'b110100_0011; next_rd = same; end
			10'b100_01011_0_0: begin code = 10'b110100_1101; next_rd = flip; end
			10'b100_01011_1_0: begin code = 10'b110100_0010; next_rd = flip; end
			10'b101_01011_0_0: begin code = 10'b110100_1010; next_rd = same; end
			10'b101_01011_1_0: begin code = 10'b110100_1010; next_rd = same; end
			10'b110_01011_0_0: begin code = 10'b110100_0110; next_rd = same; end
			10'b110_01011_1_0: begin code = 10'b110100_0110; next_rd = same; end
			10'b111_01011_0_0: begin code = 10'b110100_1110; next_rd = flip; end
			10'b111_01011_1_0: begin code = 10'b110100_1000; next_rd = flip; end
			10'b000_10000_0_0: begin code = 10'b011011_0100; next_rd = same; end
			10'b000_10000_1_0: begin code = 10'b100100_1011; next_rd = same; end
			10'b001_10000_0_0: begin code = 10'b011011_1001; next_rd = flip; end
			10'b001_10000_1_0: begin code = 10'b100100_1001; next_rd = flip; end
			10'b010_10000_0_0: begin code = 10'b011011_0101; next_rd = flip; end
			10'b010_10000_1_0: begin code = 10'b100100_0101; next_rd = flip; end
			10'b011_10000_0_0: begin code = 10'b011011_0011; next_rd = flip; end
			10'b011_10000_1_0: begin code = 10'b100100_1100; next_rd = flip; end
			10'b100_10000_0_0: begin code = 10'b011011_0010; next_rd = same; end
			10'b100_10000_1_0: begin code = 10'b100100_1101; next_rd = same; end
			10'b101_10000_0_0: begin code = 10'b011011_1010; next_rd = flip; end
			10'b101_10000_1_0: begin code = 10'b100100_1010; next_rd = flip; end
			10'b110_10000_0_0: begin code = 10'b011011_0110; next_rd = flip; end
			10'b110_10000_1_0: begin code = 10'b100100_0110; next_rd = flip; end
			10'b111_10000_0_0: begin code = 10'b011011_0001; next_rd = same; end
			10'b111_10000_1_0: begin code = 10'b100100_1110; next_rd = same; end
			10'b000_10001_0_0: begin code = 10'b100011_1011; next_rd = flip; end
			10'b000_10001_1_0: begin code = 10'b100011_0100; next_rd = flip; end
			10'b001_10001_0_0: begin code = 10'b100011_1001; next_rd = same; end
			10'b001_10001_1_0: begin code = 10'b100011_1001; next_rd = same; end
			10'b010_10001_0_0: begin code = 10'b100011_0101; next_rd = same; end
			10'b010_10001_1_0: begin code = 10'b100011_0101; next_rd = same; end
			10'b011_10001_0_0: begin code = 10'b100011_1100; next_rd = same; end
			10'b011_10001_1_0: begin code = 10'b100011_0011; next_rd = same; end
			10'b100_10001_0_0: begin code = 10'b100011_1101; next_rd = flip; end
			10'b100_10001_1_0: begin code = 10'b100011_0010; next_rd = flip; end
			10'b101_10001_0_0: begin code = 10'b100011_1010; next_rd = same; end
			10'b101_10001_1_0: begin code = 10'b100011_1010; next_rd = same; end
			10'b110_10001_0_0: begin code = 10'b100011_0110; next_rd = same; end
			10'b110_10001_1_0: begin code = 10'b100011_0110; next_rd = same; end
			10'b111_10001_0_0: begin code = 10'b100011_0111; next_rd = flip; end
			10'b111_10001_1_0: begin code = 10'b100011_0001; next_rd = flip; end
			10'b000_10010_0_0: begin code = 10'b010011_1011; next_rd = flip; end
			10'b000_10010_1_0: begin code = 10'b010011_0100; next_rd = flip; end
			10'b001_10010_0_0: begin code = 10'b010011_1001; next_rd = same; end
			10'b001_10010_1_0: begin code = 10'b010011_1001; next_rd = same; end
			10'b010_10010_0_0: begin code = 10'b010011_0101; next_rd = same; end
			10'b010_10010_1_0: begin code = 10'b010011_0101; next_rd = same; end
			10'b011_10010_0_0: begin code = 10'b010011_1100; next_rd = same; end
			10'b011_10010_1_0: begin code = 10'b010011_0011; next_rd = same; end
			10'b100_10010_0_0: begin code = 10'b010011_1101; next_rd = flip; end
			10'b100_10010_1_0: begin code = 10'b010011_0010; next_rd = flip; end
			10'b101_10010_0_0: begin code = 10'b010011_1010; next_rd = same; end
			10'b101_10010_1_0: begin code = 10'b010011_1010; next_rd = same; end
			10'b110_10010_0_0: begin code = 10'b010011_0110; next_rd = same; end
			10'b110_10010_1_0: begin code = 10'b010011_0110; next_rd = same; end
			10'b111_10010_0_0: begin code = 10'b010011_0111; next_rd = flip; end
			10'b111_10010_1_0: begin code = 10'b010011_0001; next_rd = flip; end
			10'b000_10011_0_0: begin code = 10'b110010_1011; next_rd = flip; end
			10'b000_10011_1_0: begin code = 10'b110010_0100; next_rd = flip; end
			10'b001_10011_0_0: begin code = 10'b110010_1001; next_rd = same; end
			10'b001_10011_1_0: begin code = 10'b110010_1001; next_rd = same; end
			10'b010_10011_0_0: begin code = 10'b110010_0101; next_rd = same; end
			10'b010_10011_1_0: begin code = 10'b110010_0101; next_rd = same; end
			10'b011_10011_0_0: begin code = 10'b110010_1100; next_rd = same; end
			10'b011_10011_1_0: begin code = 10'b110010_0011; next_rd = same; end
			10'b100_10011_0_0: begin code = 10'b110010_1101; next_rd = flip; end
			10'b100_10011_1_0: begin code = 10'b110010_0010; next_rd = flip; end
			10'b101_10011_0_0: begin code = 10'b110010_1010; next_rd = same; end
			10'b101_10011_1_0: begin code = 10'b110010_1010; next_rd = same; end
			10'b110_10011_0_0: begin code = 10'b110010_0110; next_rd = same; end
			10'b110_10011_1_0: begin code = 10'b110010_0110; next_rd = same; end
			10'b111_10011_0_0: begin code = 10'b110010_1110; next_rd = flip; end
			10'b111_10011_1_0: begin code = 10'b110010_0001; next_rd = flip; end
			10'b000_11000_0_0: begin code = 10'b110011_0100; next_rd = same; end
			10'b000_11000_1_0: begin code = 10'b001100_1011; next_rd = same; end
			10'b001_11000_0_0: begin code = 10'b110011_1001; next_rd = flip; end
			10'b001_11000_1_0: begin code = 10'b001100_1001; next_rd = flip; end
			10'b010_11000_0_0: begin code = 10'b110011_0101; next_rd = flip; end
			10'b010_11000_1_0: begin code = 10'b001100_0101; next_rd = flip; end
			10'b011_11000_0_0: begin code = 10'b110011_0011; next_rd = flip; end
			10'b011_11000_1_0: begin code = 10'b001100_1100; next_rd = flip; end
			10'b100_11000_0_0: begin code = 10'b110011_0010; next_rd = same; end
			10'b100_11000_1_0: begin code = 10'b001100_1101; next_rd = same; end
			10'b101_11000_0_0: begin code = 10'b110011_1010; next_rd = flip; end
			10'b101_11000_1_0: begin code = 10'b001100_1010; next_rd = flip; end
			10'b110_11000_0_0: begin code = 10'b110011_0110; next_rd = flip; end
			10'b110_11000_1_0: begin code = 10'b001100_0110; next_rd = flip; end
			10'b111_11000_0_0: begin code = 10'b110011_0001; next_rd = same; end
			10'b111_11000_1_0: begin code = 10'b001100_1110; next_rd = same; end
			10'b000_11001_0_0: begin code = 10'b100110_1011; next_rd = flip; end
			10'b000_11001_1_0: begin code = 10'b100110_0100; next_rd = flip; end
			10'b001_11001_0_0: begin code = 10'b100110_1001; next_rd = same; end
			10'b001_11001_1_0: begin code = 10'b100110_1001; next_rd = same; end
			10'b010_11001_0_0: begin code = 10'b100110_0101; next_rd = same; end
			10'b010_11001_1_0: begin code = 10'b100110_0101; next_rd = same; end
			10'b011_11001_0_0: begin code = 10'b100110_1100; next_rd = same; end
			10'b011_11001_1_0: begin code = 10'b100110_0011; next_rd = same; end
			10'b100_11001_0_0: begin code = 10'b100110_1101; next_rd = flip; end
			10'b100_11001_1_0: begin code = 10'b100110_0010; next_rd = flip; end
			10'b101_11001_0_0: begin code = 10'b100110_1010; next_rd = same; end
			10'b101_11001_1_0: begin code = 10'b100110_1010; next_rd = same; end
			10'b110_11001_0_0: begin code = 10'b100110_0110; next_rd = same; end
			10'b110_11001_1_0: begin code = 10'b100110_0110; next_rd = same; end
			10'b111_11001_0_0: begin code = 10'b100110_1110; next_rd = flip; end
			10'b111_11001_1_0: begin code = 10'b100110_0001; next_rd = flip; end
			10'b000_11010_0_0: begin code = 10'b010110_1011; next_rd = flip; end
			10'b000_11010_1_0: begin code = 10'b010110_0100; next_rd = flip; end
			10'b001_11010_0_0: begin code = 10'b010110_1001; next_rd = same; end
			10'b001_11010_1_0: begin code = 10'b010110_1001; next_rd = same; end
			10'b010_11010_0_0: begin code = 10'b010110_0101; next_rd = same; end
			10'b010_11010_1_0: begin code = 10'b010110_0101; next_rd = same; end
			10'b011_11010_0_0: begin code = 10'b010110_1100; next_rd = same; end
			10'b011_11010_1_0: begin code = 10'b010110_0011; next_rd = same; end
			10'b100_11010_0_0: begin code = 10'b010110_1101; next_rd = flip; end
			10'b100_11010_1_0: begin code = 10'b010110_0010; next_rd = flip; end
			10'b101_11010_0_0: begin code = 10'b010110_1010; next_rd = same; end
			10'b101_11010_1_0: begin code = 10'b010110_1010; next_rd = same; end
			10'b110_11010_0_0: begin code = 10'b010110_0110; next_rd = same; end
			10'b110_11010_1_0: begin code = 10'b010110_0110; next_rd = same; end
			10'b111_11010_0_0: begin code = 10'b010110_1110; next_rd = flip; end
			10'b111_11010_1_0: begin code = 10'b010110_0001; next_rd = flip; end
			10'b000_11011_0_0: begin code = 10'b110110_0100; next_rd = same; end
			10'b000_11011_1_0: begin code = 10'b001001_1011; next_rd = same; end
			10'b001_11011_0_0: begin code = 10'b110110_1001; next_rd = flip; end
			10'b001_11011_1_0: begin code = 10'b001001_1001; next_rd = flip; end
			10'b010_11011_0_0: begin code = 10'b110110_0101; next_rd = flip; end
			10'b010_11011_1_0: begin code = 10'b001001_0101; next_rd = flip; end
			10'b011_11011_0_0: begin code = 10'b110110_0011; next_rd = flip; end
			10'b011_11011_1_0: begin code = 10'b001001_1100; next_rd = flip; end
			10'b100_11011_0_0: begin code = 10'b110110_0010; next_rd = same; end
			10'b100_11011_1_0: begin code = 10'b001001_1101; next_rd = same; end
			10'b101_11011_0_0: begin code = 10'b110110_1010; next_rd = flip; end
			10'b101_11011_1_0: begin code = 10'b001001_1010; next_rd = flip; end
			10'b110_11011_0_0: begin code = 10'b110110_0110; next_rd = flip; end
			10'b110_11011_1_0: begin code = 10'b001001_0110; next_rd = flip; end
			10'b111_11011_0_0: begin code = 10'b110110_0001; next_rd = same; end
			10'b111_11011_1_0: begin code = 10'b001001_1110; next_rd = same; end
			10'b000_01100_0_0: begin code = 10'b001101_1011; next_rd = flip; end
			10'b000_01100_1_0: begin code = 10'b001101_0100; next_rd = flip; end
			10'b001_01100_0_0: begin code = 10'b001101_1001; next_rd = same; end
			10'b001_01100_1_0: begin code = 10'b001101_1001; next_rd = same; end
			10'b010_01100_0_0: begin code = 10'b001101_0101; next_rd = same; end
			10'b010_01100_1_0: begin code = 10'b001101_0101; next_rd = same; end
			10'b011_01100_0_0: begin code = 10'b001101_1100; next_rd = same; end
			10'b011_01100_1_0: begin code = 10'b001101_0011; next_rd = same; end
			10'b100_01100_0_0: begin code = 10'b001101_1101; next_rd = flip; end
			10'b100_01100_1_0: begin code = 10'b001101_0010; next_rd = flip; end
			10'b101_01100_0_0: begin code = 10'b001101_1010; next_rd = same; end
			10'b101_01100_1_0: begin code = 10'b001101_1010; next_rd = same; end
			10'b110_01100_0_0: begin code = 10'b001101_0110; next_rd = same; end
			10'b110_01100_1_0: begin code = 10'b001101_0110; next_rd = same; end
			10'b111_01100_0_0: begin code = 10'b001101_1110; next_rd = flip; end
			10'b111_01100_1_0: begin code = 10'b001101_0001; next_rd = flip; end
			10'b000_01101_0_0: begin code = 10'b101100_1011; next_rd = flip; end
			10'b000_01101_1_0: begin code = 10'b101100_0100; next_rd = flip; end
			10'b001_01101_0_0: begin code = 10'b101100_1001; next_rd = same; end
			10'b001_01101_1_0: begin code = 10'b101100_1001; next_rd = same; end
			10'b010_01101_0_0: begin code = 10'b101100_0101; next_rd = same; end
			10'b010_01101_1_0: begin code = 10'b101100_0101; next_rd = same; end
			10'b011_01101_0_0: begin code = 10'b101100_1100; next_rd = same; end
			10'b011_01101_1_0: begin code = 10'b101100_0011; next_rd = same; end
			10'b100_01101_0_0: begin code = 10'b101100_1101; next_rd = flip; end
			10'b100_01101_1_0: begin code = 10'b101100_0010; next_rd = flip; end
			10'b101_01101_0_0: begin code = 10'b101100_1010; next_rd = same; end
			10'b101_01101_1_0: begin code = 10'b101100_1010; next_rd = same; end
			10'b110_01101_0_0: begin code = 10'b101100_0110; next_rd = same; end
			10'b110_01101_1_0: begin code = 10'b101100_0110; next_rd = same; end
			10'b111_01101_0_0: begin code = 10'b101100_1110; next_rd = flip; end
			10'b111_01101_1_0: begin code = 10'b101100_1000; next_rd = flip; end
			10'b000_01110_0_0: begin code = 10'b011100_1011; next_rd = flip; end
			10'b000_01110_1_0: begin code = 10'b011100_0100; next_rd = flip; end
			10'b001_01110_0_0: begin code = 10'b011100_1001; next_rd = same; end
			10'b001_01110_1_0: begin code = 10'b011100_1001; next_rd = same; end
			10'b010_01110_0_0: begin code = 10'b011100_0101; next_rd = same; end
			10'b010_01110_1_0: begin code = 10'b011100_0101; next_rd = same; end
			10'b011_01110_0_0: begin code = 10'b011100_1100; next_rd = same; end
			10'b011_01110_1_0: begin code = 10'b011100_0011; next_rd = same; end
			10'b100_01110_0_0: begin code = 10'b011100_1101; next_rd = flip; end
			10'b100_01110_1_0: begin code = 10'b011100_0010; next_rd = flip; end
			10'b101_01110_0_0: begin code = 10'b011100_1010; next_rd = same; end
			10'b101_01110_1_0: begin code = 10'b011100_1010; next_rd = same; end
			10'b110_01110_0_0: begin code = 10'b011100_0110; next_rd = same; end
			10'b110_01110_1_0: begin code = 10'b011100_0110; next_rd = same; end
			10'b111_01110_0_0: begin code = 10'b011100_1110; next_rd = flip; end
			10'b111_01110_1_0: begin code = 10'b011100_1000; next_rd = flip; end
			10'b000_01111_0_0: begin code = 10'b010111_0100; next_rd = same; end
			10'b000_01111_1_0: begin code = 10'b101000_1011; next_rd = same; end
			10'b001_01111_0_0: begin code = 10'b010111_1001; next_rd = flip; end
			10'b001_01111_1_0: begin code = 10'b101000_1001; next_rd = flip; end
			10'b010_01111_0_0: begin code = 10'b010111_0101; next_rd = flip; end
			10'b010_01111_1_0: begin code = 10'b101000_0101; next_rd = flip; end
			10'b011_01111_0_0: begin code = 10'b010111_0011; next_rd = flip; end
			10'b011_01111_1_0: begin code = 10'b101000_1100; next_rd = flip; end
			10'b100_01111_0_0: begin code = 10'b010111_0010; next_rd = same; end
			10'b100_01111_1_0: begin code = 10'b101000_1101; next_rd = same; end
			10'b101_01111_0_0: begin code = 10'b010111_1010; next_rd = flip; end
			10'b101_01111_1_0: begin code = 10'b101000_1010; next_rd = flip; end
			10'b110_01111_0_0: begin code = 10'b010111_0110; next_rd = flip; end
			10'b110_01111_1_0: begin code = 10'b101000_0110; next_rd = flip; end
			10'b111_01111_0_0: begin code = 10'b010111_0001; next_rd = same; end
			10'b111_01111_1_0: begin code = 10'b101000_1110; next_rd = same; end
			10'b000_10100_0_0: begin code = 10'b001011_1011; next_rd = flip; end
			10'b000_10100_1_0: begin code = 10'b001011_0100; next_rd = flip; end
			10'b001_10100_0_0: begin code = 10'b001011_1001; next_rd = same; end
			10'b001_10100_1_0: begin code = 10'b001011_1001; next_rd = same; end
			10'b010_10100_0_0: begin code = 10'b001011_0101; next_rd = same; end
			10'b010_10100_1_0: begin code = 10'b001011_0101; next_rd = same; end
			10'b011_10100_0_0: begin code = 10'b001011_1100; next_rd = same; end
			10'b011_10100_1_0: begin code = 10'b001011_0011; next_rd = same; end
			10'b100_10100_0_0: begin code = 10'b001011_1101; next_rd = flip; end
			10'b100_10100_1_0: begin code = 10'b001011_0010; next_rd = flip; end
			10'b101_10100_0_0: begin code = 10'b001011_1010; next_rd = same; end
			10'b101_10100_1_0: begin code = 10'b001011_1010; next_rd = same; end
			10'b110_10100_0_0: begin code = 10'b001011_0110; next_rd = same; end
			10'b110_10100_1_0: begin code = 10'b001011_0110; next_rd = same; end
			10'b111_10100_0_0: begin code = 10'b001011_0111; next_rd = flip; end
			10'b111_10100_1_0: begin code = 10'b001011_0001; next_rd = flip; end
			10'b000_10101_0_0: begin code = 10'b101010_1011; next_rd = flip; end
			10'b000_10101_1_0: begin code = 10'b101010_0100; next_rd = flip; end
			10'b001_10101_0_0: begin code = 10'b101010_1001; next_rd = same; end
			10'b001_10101_1_0: begin code = 10'b101010_1001; next_rd = same; end
			10'b010_10101_0_0: begin code = 10'b101010_0101; next_rd = same; end
			10'b010_10101_1_0: begin code = 10'b101010_0101; next_rd = same; end
			10'b011_10101_0_0: begin code = 10'b101010_1100; next_rd = same; end
			10'b011_10101_1_0: begin code = 10'b101010_0011; next_rd = same; end
			10'b100_10101_0_0: begin code = 10'b101010_1101; next_rd = flip; end
			10'b100_10101_1_0: begin code = 10'b101010_0010; next_rd = flip; end
			10'b101_10101_0_0: begin code = 10'b101010_1010; next_rd = same; end
			10'b101_10101_1_0: begin code = 10'b101010_1010; next_rd = same; end
			10'b110_10101_0_0: begin code = 10'b101010_0110; next_rd = same; end
			10'b110_10101_1_0: begin code = 10'b101010_0110; next_rd = same; end
			10'b111_10101_0_0: begin code = 10'b101010_1110; next_rd = flip; end
			10'b111_10101_1_0: begin code = 10'b101010_0001; next_rd = flip; end
			10'b000_10110_0_0: begin code = 10'b011010_1011; next_rd = flip; end
			10'b000_10110_1_0: begin code = 10'b011010_0100; next_rd = flip; end
			10'b001_10110_0_0: begin code = 10'b011010_1001; next_rd = same; end
			10'b001_10110_1_0: begin code = 10'b011010_1001; next_rd = same; end
			10'b010_10110_0_0: begin code = 10'b011010_0101; next_rd = same; end
			10'b010_10110_1_0: begin code = 10'b011010_0101; next_rd = same; end
			10'b011_10110_0_0: begin code = 10'b011010_1100; next_rd = same; end
			10'b011_10110_1_0: begin code = 10'b011010_0011; next_rd = same; end
			10'b100_10110_0_0: begin code = 10'b011010_1101; next_rd = flip; end
			10'b100_10110_1_0: begin code = 10'b011010_0010; next_rd = flip; end
			10'b101_10110_0_0: begin code = 10'b011010_1010; next_rd = same; end
			10'b101_10110_1_0: begin code = 10'b011010_1010; next_rd = same; end
			10'b110_10110_0_0: begin code = 10'b011010_0110; next_rd = same; end
			10'b110_10110_1_0: begin code = 10'b011010_0110; next_rd = same; end
			10'b111_10110_0_0: begin code = 10'b011010_1110; next_rd = flip; end
			10'b111_10110_1_0: begin code = 10'b011010_0001; next_rd = flip; end
			10'b000_10111_0_0: begin code = 10'b111010_0100; next_rd = same; end
			10'b000_10111_1_0: begin code = 10'b000101_1011; next_rd = same; end
			10'b001_10111_0_0: begin code = 10'b111010_1001; next_rd = flip; end
			10'b001_10111_1_0: begin code = 10'b000101_1001; next_rd = flip; end
			10'b010_10111_0_0: begin code = 10'b111010_0101; next_rd = flip; end
			10'b010_10111_1_0: begin code = 10'b000101_0101; next_rd = flip; end
			10'b011_10111_0_0: begin code = 10'b111010_0011; next_rd = flip; end
			10'b011_10111_1_0: begin code = 10'b000101_1100; next_rd = flip; end
			10'b100_10111_0_0: begin code = 10'b111010_0010; next_rd = same; end
			10'b100_10111_1_0: begin code = 10'b000101_1101; next_rd = same; end
			10'b101_10111_0_0: begin code = 10'b111010_1010; next_rd = flip; end
			10'b101_10111_1_0: begin code = 10'b000101_1010; next_rd = flip; end
			10'b110_10111_0_0: begin code = 10'b111010_0110; next_rd = flip; end
			10'b110_10111_1_0: begin code = 10'b000101_0110; next_rd = flip; end
			10'b111_10111_0_0: begin code = 10'b111010_0001; next_rd = same; end
			10'b111_10111_1_0: begin code = 10'b000101_1110; next_rd = same; end
			10'b000_11100_0_0: begin code = 10'b001110_1011; next_rd = flip; end
			10'b000_11100_1_0: begin code = 10'b001110_0100; next_rd = flip; end
			10'b001_11100_0_0: begin code = 10'b001110_1001; next_rd = same; end
			10'b001_11100_1_0: begin code = 10'b001110_1001; next_rd = same; end
			10'b010_11100_0_0: begin code = 10'b001110_0101; next_rd = same; end
			10'b010_11100_1_0: begin code = 10'b001110_0101; next_rd = same; end
			10'b011_11100_0_0: begin code = 10'b001110_1100; next_rd = same; end
			10'b011_11100_1_0: begin code = 10'b001110_0011; next_rd = same; end
			10'b100_11100_0_0: begin code = 10'b001110_1101; next_rd = flip; end
			10'b100_11100_1_0: begin code = 10'b001110_0010; next_rd = flip; end
			10'b101_11100_0_0: begin code = 10'b001110_1010; next_rd = same; end
			10'b101_11100_1_0: begin code = 10'b001110_1010; next_rd = same; end
			10'b110_11100_0_0: begin code = 10'b001110_0110; next_rd = same; end
			10'b110_11100_1_0: begin code = 10'b001110_0110; next_rd = same; end
			10'b111_11100_0_0: begin code = 10'b001110_1110; next_rd = flip; end
			10'b111_11100_1_0: begin code = 10'b001110_0001; next_rd = flip; end
			10'b000_11101_0_0: begin code = 10'b101110_0100; next_rd = same; end
			10'b000_11101_1_0: begin code = 10'b010001_1011; next_rd = same; end
			10'b001_11101_0_0: begin code = 10'b101110_1001; next_rd = flip; end
			10'b001_11101_1_0: begin code = 10'b010001_1001; next_rd = flip; end
			10'b010_11101_0_0: begin code = 10'b101110_0101; next_rd = flip; end
			10'b010_11101_1_0: begin code = 10'b010001_0101; next_rd = flip; end
			10'b011_11101_0_0: begin code = 10'b101110_0011; next_rd = flip; end
			10'b011_11101_1_0: begin code = 10'b010001_1100; next_rd = flip; end
			10'b100_11101_0_0: begin code = 10'b101110_0010; next_rd = same; end
			10'b100_11101_1_0: begin code = 10'b010001_1101; next_rd = same; end
			10'b101_11101_0_0: begin code = 10'b101110_1010; next_rd = flip; end
			10'b101_11101_1_0: begin code = 10'b010001_1010; next_rd = flip; end
			10'b110_11101_0_0: begin code = 10'b101110_0110; next_rd = flip; end
			10'b110_11101_1_0: begin code = 10'b010001_0110; next_rd = flip; end
			10'b111_11101_0_0: begin code = 10'b101110_0001; next_rd = same; end
			10'b111_11101_1_0: begin code = 10'b010001_1110; next_rd = same; end
			10'b000_11110_0_0: begin code = 10'b011110_0100; next_rd = same; end
			10'b000_11110_1_0: begin code = 10'b100001_1011; next_rd = same; end
			10'b001_11110_0_0: begin code = 10'b011110_1001; next_rd = flip; end
			10'b001_11110_1_0: begin code = 10'b100001_1001; next_rd = flip; end
			10'b010_11110_0_0: begin code = 10'b011110_0101; next_rd = flip; end
			10'b010_11110_1_0: begin code = 10'b100001_0101; next_rd = flip; end
			10'b011_11110_0_0: begin code = 10'b011110_0011; next_rd = flip; end
			10'b011_11110_1_0: begin code = 10'b100001_1100; next_rd = flip; end
			10'b100_11110_0_0: begin code = 10'b011110_0010; next_rd = same; end
			10'b100_11110_1_0: begin code = 10'b100001_1101; next_rd = same; end
			10'b101_11110_0_0: begin code = 10'b011110_1010; next_rd = flip; end
			10'b101_11110_1_0: begin code = 10'b100001_1010; next_rd = flip; end
			10'b110_11110_0_0: begin code = 10'b011110_0110; next_rd = flip; end
			10'b110_11110_1_0: begin code = 10'b100001_0110; next_rd = flip; end
			10'b111_11110_0_0: begin code = 10'b011110_0001; next_rd = same; end
			10'b111_11110_1_0: begin code = 10'b100001_1110; next_rd = same; end
			10'b000_11111_0_0: begin code = 10'b101011_0100; next_rd = same; end
			10'b000_11111_1_0: begin code = 10'b010100_1011; next_rd = same; end
			10'b001_11111_0_0: begin code = 10'b101011_1001; next_rd = flip; end
			10'b001_11111_1_0: begin code = 10'b010100_1001; next_rd = flip; end
			10'b010_11111_0_0: begin code = 10'b101011_0101; next_rd = flip; end
			10'b010_11111_1_0: begin code = 10'b010100_0101; next_rd = flip; end
			10'b011_11111_0_0: begin code = 10'b101011_0011; next_rd = flip; end
			10'b011_11111_1_0: begin code = 10'b010100_1100; next_rd = flip; end
			10'b100_11111_0_0: begin code = 10'b101011_0010; next_rd = same; end
			10'b100_11111_1_0: begin code = 10'b010100_1101; next_rd = same; end
			10'b101_11111_0_0: begin code = 10'b101011_1010; next_rd = flip; end
			10'b101_11111_1_0: begin code = 10'b010100_1010; next_rd = flip; end
			10'b110_11111_0_0: begin code = 10'b101011_0110; next_rd = flip; end
			10'b110_11111_1_0: begin code = 10'b010100_0110; next_rd = flip; end
			10'b111_11111_0_0: begin code = 10'b101011_0001; next_rd = same; end
			10'b111_11111_1_0: begin code = 10'b010100_1110; next_rd = same; end
					
			10'b000_11100_0_1: begin code = 10'b001111_0100; next_rd = same; end
			10'b000_11100_1_1: begin code = 10'b110000_1011; next_rd = same; end
			10'b001_11100_0_1: begin code = 10'b001111_1001; next_rd = flip; end
			10'b001_11100_1_1: begin code = 10'b110000_0110; next_rd = flip; end
			10'b010_11100_0_1: begin code = 10'b001111_0101; next_rd = flip; end
			10'b010_11100_1_1: begin code = 10'b110000_1010; next_rd = flip; end
			10'b011_11100_0_1: begin code = 10'b001111_0011; next_rd = flip; end
			10'b011_11100_1_1: begin code = 10'b110000_1100; next_rd = flip; end
			10'b100_11100_0_1: begin code = 10'b001111_0010; next_rd = same; end
			10'b100_11100_1_1: begin code = 10'b110000_1101; next_rd = same; end
			10'b101_11100_0_1: begin code = 10'b001111_1010; next_rd = flip; end
			10'b101_11100_1_1: begin code = 10'b110000_0101; next_rd = flip; end
			10'b110_11100_0_1: begin code = 10'b001111_0110; next_rd = flip; end
			10'b110_11100_1_1: begin code = 10'b110000_1001; next_rd = flip; end
			10'b111_11100_0_1: begin code = 10'b001111_1000; next_rd = same; end
			10'b111_11100_1_1: begin code = 10'b110000_0111; next_rd = same; end
			10'b111_10111_0_1: begin code = 10'b111010_1000; next_rd = same; end
			10'b111_10111_1_1: begin code = 10'b000101_0111; next_rd = same; end
			10'b111_11011_0_1: begin code = 10'b110110_1000; next_rd = same; end
			10'b111_11011_1_1: begin code = 10'b001001_0111; next_rd = same; end
			10'b111_11101_0_1: begin code = 10'b101110_1000; next_rd = same; end
			10'b111_11101_1_1: begin code = 10'b010001_0111; next_rd = same; end
			10'b111_11110_0_1: begin code = 10'b011110_1000; next_rd = same; end
			10'b111_11110_1_1: begin code = 10'b100001_0111; next_rd = same; end		
			
			default: begin code = 10'b0; next_rd = same; end
		endcase
	end

endmodule
