
module clock_divider (

	input      inclk0,
	output reg clk_out

);

	parameter WIDTH = 4;

	reg [WIDTH - 1 : 0] counter = 4'b0;

	

endmodule